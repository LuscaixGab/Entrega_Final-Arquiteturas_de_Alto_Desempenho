module num #(
	parameter N = 0)(
	output [13:0] n);
	
	assign n = N;
	
endmodule